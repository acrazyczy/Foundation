`include "constant.vh"

module RS(
    input wire clk_in,
    input wire rst_in,
    input wire rdy_in,


);
endmodule : RS