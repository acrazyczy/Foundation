`include "constant.vh"

module rob(
    input clk_in,
    input rst_in,
    input rdy_in,

    
);
endmodule : rob