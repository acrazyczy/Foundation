`ifndef _constant_h
`define _constant_h
`define IDWidth 32
`define AddressWidth 32
`endif