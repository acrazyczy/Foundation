`include "constant.vh"

module lbuffer(
    input wire clk_in,
    input wire rst_in,
    input wire rdy_in,
);
endmodule : lbuffer